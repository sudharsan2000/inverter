* SPICE3 file created from inv.ext - technology: scmos

.option scale=1u

M1000 out in gnd Gnd nfet w=4 l=2
+  ad=28 pd=22 as=28 ps=22
M1001 out in vdd vdd pfet w=8 l=2
+  ad=56 pd=30 as=40 ps=26
C0 gnd Gnd 2.26fF
C1 out Gnd 2.26fF
C2 in Gnd 4.37fF
